//名称：指令译码器
//input：code(输入32位数据)
//output:instruct(32位译码后的串)

module Decoder(
    input [31:0] code,
    output reg [31:0] instruct
);
    wire [5:0] op;
    wire [5:0] func;
    assign op=code[31:26];
    assign func=code[5:0];

    always @(*) 
    begin
        case(op)
            6'b000000:
            begin
                case(func)
                    6'b100000: instruct = 32'b00000000_00000000_00000000_00000001; //add
                    6'b100001: instruct = 32'b00000000_00000000_00000000_00000010; //addu
                    6'b100010: instruct = 32'b00000000_00000000_00000000_00000100; //sub
                    6'b100011: instruct = 32'b00000000_00000000_00000000_00001000; //subu
                    6'b100100: instruct = 32'b00000000_00000000_00000000_00010000; //and
                    6'b100101: instruct = 32'b00000000_00000000_00000000_00100000; //or
                    6'b100110: instruct = 32'b00000000_00000000_00000000_01000000; //xor
                    6'b100111: instruct = 32'b00000000_00000000_00000000_10000000; //nor
                    6'b101010: instruct = 32'b00000000_00000000_00000001_00000000; //slt
                    6'b101011: instruct = 32'b00000000_00000000_00000010_00000000; //sltu
                    6'b000000: instruct = 32'b00000000_00000000_00000100_00000000; //sll
                    6'b000010: instruct = 32'b00000000_00000000_00001000_00000000; //srl
                    6'b000011: instruct = 32'b00000000_00000000_00010000_00000000; //sra
                    6'b000100: instruct = 32'b00000000_00000000_00100000_00000000; //sllv
                    6'b000110: instruct = 32'b00000000_00000000_01000000_00000000; //srlv
                    6'b000111: instruct = 32'b00000000_00000000_10000000_00000000; //srav
                    6'b001000: instruct = 32'b00000000_00000001_00000000_00000000; //jr
                    default: instruct = 32'b0;
                endcase
            end
            6'b001000: instruct = 32'b00000000_00000010_00000000_00000000; //addi
            6'b001001: instruct = 32'b00000000_00000100_00000000_00000000; //addiu
            6'b001100: instruct = 32'b00000000_00001000_00000000_00000000; //andi
            6'b001101: instruct = 32'b00000000_00010000_00000000_00000000; //ori
            6'b001110: instruct = 32'b00000000_00100000_00000000_00000000; //xori
            6'b100011: instruct = 32'b00000000_01000000_00000000_00000000; //lw
            6'b101011: instruct = 32'b00000000_10000000_00000000_00000000; //sw
            6'b000100: instruct = 32'b00000001_00000000_00000000_00000000; //beq
            6'b000101: instruct = 32'b00000010_00000000_00000000_00000000; //bne
            6'b001010: instruct = 32'b00000100_00000000_00000000_00000000; //slti
            6'b001011: instruct = 32'b00001000_00000000_00000000_00000000; //sltiu
            6'b001111: instruct = 32'b00010000_00000000_00000000_00000000; //lui
            6'b000010: instruct = 32'b00100000_00000000_00000000_00000000; //j
            6'b000011: instruct = 32'b01000000_00000000_00000000_00000000; //jal
            default: instruct = 32'b0;
        endcase
    end
endmodule